module bnot(input a, output r);
    assign r = ~a;
endmodule