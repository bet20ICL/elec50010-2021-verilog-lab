module multiplier_parallel_tb();
    logic clk;
    
    initial begin
        $dumpfile("multiplier_pipelined.vcd");
    end