module ram256x8(
    input logic clk,
    input logic write,
    input logic [7:0] addr,
    input logic [7:0] data_in,
    output logic [7:0] data_out,
)

endmodule