module opcode_decoder(
    input clk,
    input logic[5:0] opcode,
    output rtype,
    output itype,
    output jtype
);

    always_comb begin
        
    end

endmodule